module fsk_demodulator(
    input clk,           // ʱ���ź�
    input fsk_in,        // FSK��������
    output reg data_out  // �������������
);

// ��������
parameter COUNTER_MAX = 10000;  // �����������ֵ
parameter PERIODS_TO_MEASURE = 2;  // Ҫ������������
parameter THRESHOLD0 = 80 * PERIODS_TO_MEASURE;    //160 ��ֵ�������ж����ĸ�����
parameter THRESHOLD1 = 93 * PERIODS_TO_MEASURE;    //186 ��ֵ�������ж����ĸ�����
parameter THRESHOLD2 = 97;    // ��ֵ�������ж����ĸ�����
parameter THRESHOLD3 = 103;    // ��ֵ�������ж����ĸ�����
parameter PERIODS_NOISE = 10;  // ����������

// �ڲ��źŶ���
reg [13:0] counter = 0;         // �����������ڲ������ڳ���
reg fsk_in_last = 0;            // ��һ��ʱ�����ڵ�FSK����
reg [15:0] period_sum = 0;      // �����������ڳ���֮��
reg [8:0] periods_measured = 0; // �Ѳ�����������


 
 
 
initial begin
	data_out = 0;
	//clk_out = 0;
end

// ����FSK�źŵ����ڳ��Ȳ��ۼ�
always @(posedge clk) begin
    fsk_in_last <= fsk_in;
    if ((periods_measured == 0 || counter > PERIODS_NOISE)) begin
		if (periods_measured < PERIODS_TO_MEASURE) begin
			period_sum <= period_sum + counter;
			periods_measured <= periods_measured + 1;
		end
		counter <= 0;
    end else begin
        if (counter < COUNTER_MAX) begin
            counter <= counter + 1;
        end else begin
			// �����ۼ����ͼ�����
			counter = 0;
			period_sum <= 0;
			periods_measured <= 0;
        end
    end

    if (periods_measured >= PERIODS_TO_MEASURE) begin
        if (period_sum > THRESHOLD0 && period_sum < THRESHOLD1) begin
            data_out <= 1;  // ���յ�����1
        end else begin
            data_out <= 0;  // ���յ�����0
        end
        // �����ۼ����ͼ�����
        period_sum <= 0;
        periods_measured <= 0;
    end
end

endmodule
